//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU function code definiRons
// Author:  rz
// Last rev. 24/06/2024
//-----------------------------------------------------


`define RADD        2'b00
`define RMUL        2'b01
`define RDIVIDED    2'b10
`define RNOP    2'b11